// ============================================================================
// top_dsa_seq.sv  — top con Virtual JTAG, LEDs de estado y BRAMs
// ============================================================================

`timescale 1ps/1ps
`define MEM_INIT_FILE "img_in_64x64.hex"

module top_dsa_seq
#(
  parameter int AW                = 12,
  parameter int DEB_W             = 20,      // debounce (~10–20 ms @50MHz)
  parameter int RST_STRETCH_W     = 22
)(
  input  logic clk_50,
  input  logic rst_n,          // reset asíncrono activo bajo
  input  logic start_sw,       // switch físico (opcional)

  output logic led_done,       // latched hasta nuevo start/reset
  output logic led_reset_evt,  // pulso tras reset (visual)
  output logic led_start_on    // nivel del start_sw filtrado
);

  // ---------------- Señales core ----------------
  logic        start_pulse_sw;
  logic        start_pulse_jtag;
  logic        busy, done;

  logic [15:0] in_w_cfg, in_h_cfg, scale_q88_cfg; // JTAG
  logic [15:0] in_w, in_h, scale_q88;             // hacia core

  logic [15:0] out_w_s, out_h_s;

  logic [AW-1:0] in_raddr_core;
  logic [7:0]    in_rdata;

  logic [AW-1:0] out_waddr;
  logic [7:0]    out_wdata;
  logic          out_we;

  // =======================================================================
  // 1) Virtual JTAG + wrapper jtag_connect (control + lectura BRAMs)
  // =======================================================================
  // Señales del IP vJTAG
  wire tck, tdi, tdo;
  wire [1:0] ir_in, ir_out;
  wire vs_cdr, vs_sdr, vs_e1dr, vs_pdr, vs_e2dr, vs_udr, vs_cir, vs_uir;

  vjtag u_vjtag (
    .tdi                (tdi),
    .tdo                (tdo),
    .ir_in              (ir_in),
    .ir_out             (ir_out),
    .virtual_state_cdr  (vs_cdr),
    .virtual_state_sdr  (vs_sdr),
    .virtual_state_e1dr (vs_e1dr),
    .virtual_state_pdr  (vs_pdr),
    .virtual_state_e2dr (vs_e2dr),
    .virtual_state_udr  (vs_udr),
    .virtual_state_cir  (vs_cir),
    .virtual_state_uir  (vs_uir),
    .tck                (tck)
  );

  // Señales JTAG para lectura de BRAMs
  logic [AW-1:0] jtag_in_raddr;
  logic  [7:0]   jtag_in_rdata;
  logic [AW-1:0] jtag_out_raddr;
  logic  [7:0]   jtag_out_rdata;

  jtag_connect #(.DRW(40), .AW(AW)) u_jc (
    .tck         (tck),
    .tdi         (tdi),
    .tdo         (tdo),
    .ir_in       (ir_in),
    .ir_out      (ir_out),
    .vs_cdr      (vs_cdr),
    .vs_sdr      (vs_sdr),
    .vs_udr      (vs_udr),

    .start_pulse     (start_pulse_jtag),
    .cfg_in_w        (in_w_cfg),
    .cfg_in_h        (in_h_cfg),
    .cfg_scale_q88   (scale_q88_cfg),
    .status_done     (done),

    .in_mem_raddr    (jtag_in_raddr),
    .in_mem_rdata    (jtag_in_rdata),

    .out_mem_raddr   (jtag_out_raddr),
    .out_mem_rdata   (jtag_out_rdata),

    .clk_sys     (clk_50),
    .rst_sys_n   (rst_n)
  );

  // =========================================================================
  // 2) Sincronizador + antirrebote del switch de start
  // =========================================================================
  logic sw_meta, sw_sync;
  always_ff @(posedge clk_50 or negedge rst_n) begin
    if (!rst_n) begin
      sw_meta <= 1'b0;
      sw_sync <= 1'b0;
    end else begin
      sw_meta <= start_sw;
      sw_sync <= sw_meta;
    end
  end

  logic [DEB_W-1:0] deb_cnt;
  logic             sw_debounced, sw_debounced_q;

  always_ff @(posedge clk_50 or negedge rst_n) begin
    if (!rst_n) begin
      deb_cnt        <= '0;
      sw_debounced   <= 1'b0;
      sw_debounced_q <= 1'b0;
    end else begin
      if (sw_sync != sw_debounced) begin
        deb_cnt <= '0;
      end else if (deb_cnt != {DEB_W{1'b1}}) begin
        deb_cnt <= deb_cnt + 1'b1;
      end
      if (deb_cnt == {DEB_W{1'b1}}) begin
        sw_debounced <= sw_sync;
      end
      sw_debounced_q <= sw_debounced;
    end
  end

  assign start_pulse_sw = (sw_debounced & ~sw_debounced_q);
  assign led_start_on   = sw_debounced;

  // =========================================================================
  // 3) LED de evento de reset (latido corto)
  // =========================================================================
  logic [RST_STRETCH_W-1:0] rst_cnt;
  always_ff @(posedge clk_50 or negedge rst_n) begin
    if (!rst_n) begin
      rst_cnt <= {RST_STRETCH_W{1'b1}};
    end else begin
      if (rst_cnt != '0) rst_cnt <= rst_cnt - 1'b1;
    end
  end
  assign led_reset_evt = (rst_cnt != '0);

  // =========================================================================
  // 4) Memorias on-chip
  // =========================================================================
  // ENTRADA para el núcleo (lectura por core)
  onchip_mem_img #(
    .ADDR_W (AW),
    .INIT_EN(1'b1)
  ) mem_in (
    .clk   (clk_50),
    .raddr (in_raddr_core),
    .rdata (in_rdata),
    .waddr ('0),
    .wdata ('0),
    .we    (1'b0)
  );

  // ENTRADA "espejo" solo-lectura para JTAG (misma inicialización)
  onchip_mem_img #(
    .ADDR_W (AW),
    .INIT_EN(1'b1)
  ) mem_in_view (
    .clk   (clk_50),
    .raddr (jtag_in_raddr),
    .rdata (jtag_in_rdata),
    .waddr ('0),
    .wdata ('0),
    .we    (1'b0)
  );

  // SALIDA: escritura desde el core; lectura por JTAG
  onchip_mem_img #(
    .ADDR_W (AW),
    .INIT_EN(1'b0)
  ) mem_out (
    .clk   (clk_50),
    .raddr (jtag_out_raddr),
    .rdata (jtag_out_rdata),
    .waddr (out_waddr),
    .wdata (out_wdata),
    .we    (out_we)
  );

  // =========================================================================
  // 5) Parámetros desde JTAG
  // =========================================================================
  assign in_w      = in_w_cfg;
  assign in_h      = in_h_cfg;
  assign scale_q88 = scale_q88_cfg;

  // Start por JTAG o por switch
  wire start_any = start_pulse_jtag | start_pulse_sw;

  // =========================================================================
  // 6) Núcleo bilineal
  // =========================================================================
  bilinear_seq #(.AW(AW)) core (
    .clk         (clk_50),
    .rst_n       (rst_n),
    .start       (start_any),
    .busy        (busy),
    .done        (done),

    .i_in_w      (in_w),
    .i_in_h      (in_h),
    .i_scale_q88 (scale_q88),

    .o_out_w     (out_w_s),
    .o_out_h     (out_h_s),

    .in_raddr    (in_raddr_core),
    .in_rdata    (in_rdata),

    .out_waddr   (out_waddr),
    .out_wdata   (out_wdata),
    .out_we      (out_we)
  );

  // =========================================================================
  // 7) LED done latcheado
  // =========================================================================
  always_ff @(posedge clk_50 or negedge rst_n) begin
    if (!rst_n) begin
      led_done <= 1'b0;
    end else begin
      if (start_any)
        led_done <= 1'b0;
      else if (done)
        led_done <= 1'b1;
    end
  end

endmodule
